`ifndef DLA_DMA_PARAM_SVH
`define DLA_DMA_PARAM_SVH
  localparam string DEVICE = "AGX5";
  localparam int C_CSR_AXI_ADDR_WIDTH = 11;
  localparam int C_CSR_AXI_DATA_WIDTH = 32;
  localparam int C_DDR_AXI_ADDR_WIDTH = 32;
  localparam int C_DDR_AXI_BURST_WIDTH = 4;
  localparam int C_DDR_AXI_DATA_WIDTH = 512;
  localparam int C_DDR_AXI_THREAD_ID_WIDTH = 2;
  localparam int CONFIG_DATA_BYTES = 4;
  localparam int CONFIG_READER_DATA_BYTES = 8;
  localparam int FILTER_READER_DATA_BYTES = 64;
  localparam int FEATURE_READER_DATA_BYTES = 8;
  localparam int FEATURE_WRITER_DATA_BYTES = 8;
  localparam int CONFIG_NUM_MODULES = 16;
  localparam int MODULE_ID_WIDTH = 8;
  localparam int CONFIG_CHANNEL_WIDTH = 32;
  localparam int CONFIG_CACHE_DEPTH = 641;
  localparam int CONFIG_NETWORK_QUANTIZE_DEPTHS [255:0] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,512,64,32};
  localparam bit CONFIG_NETWORK_CROSS_CLOCK [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,1,0,0,0,0,0,1};
  localparam bit CONFIG_NETWORK_CROSS_CLOCK_AXI [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
  localparam int CONFIG_NETWORK_FIFO_MIN_DEPTH [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256};
  localparam int CONFIG_NETWORK_NUM_PIPELINE_STAGES [255:1] = {0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1};
  localparam int CONFIG_ID_PADDING = 0;
  localparam int CONFIG_ID_FILTER_READER = 1;
  localparam int CONFIG_ID_INPUT_FEEDER_MUX = 2;
  localparam int CONFIG_ID_INPUT_FEEDER_WRITER = 3;
  localparam int CONFIG_ID_INPUT_FEEDER_IN = 4;
  localparam int CONFIG_ID_INPUT_FEEDER_READER = 5;
  localparam int CONFIG_ID_INPUT_FEEDER_OUT = 6;
  localparam int CONFIG_ID_FEATURE_WRITER = 7;
  localparam int CONFIG_ID_FEATURE_READER = 8;
  localparam int CONFIG_ID_XBAR = 9;
  localparam int CONFIG_ID_ACTIVATION = 10;
  localparam int CONFIG_ID_POOL = 11;
  localparam int CONFIG_ID_SOFTMAX = 12;
  localparam int CONFIG_ID_OUTPUT_STREAMER = 13;
  localparam int CONFIG_ID_OUTPUT_STREAMER_FLUSH = 14;
  localparam int CONFIG_ID_WRITER_STREAMER_SEL = 15;
  localparam int CONFIG_ID_LAYOUT_TRANSFORM = 16;
  localparam bit ENABLE_DEBUG = 0;
  localparam bit ENABLE_INPUT_STREAMING = 1;
  localparam int AXI_ISTREAM_DATA_WIDTH = 128;
  localparam int AXI_ISTREAM_FIFO_DEPTH = 128;
  localparam bit ENABLE_ON_CHIP_PARAMETERS = 1;
  localparam bit ENABLE_MIXED_PRECISION = 0;
  localparam int KVEC_OVER_CVEC = 1;
  localparam int SB_ADDR_WIDTH = 11;
  localparam int STREAM_BUFFER_DEPTH = 2048;
  localparam bit[927:0] PE_ARRAY_PARAM_BITS = 928'h000000010000000200000001000000020000000700000007000000050000000f000000050000000f000000040000000c0000000000000001000000010000000000000001000000000000000c00000001000000010000000c00000004000000040000000000000001000000010000000100000004;
  localparam int PE_ARRAY_EXIT_FIFO_DEPTH = 512;
  localparam int SCRATCHPAD_FILTER_DEPTH = 1532;
  localparam int SCRATCHPAD_BIAS_SCALE_DEPTH = 26;
  localparam int SCRATCHPAD_NUM_FILTER_PORTS = 4;
  localparam int SCRATCHPAD_NUM_BIAS_SCALE_PORTS = 4;
  localparam int SCRATCHPAD_MEGABLOCK_WIDTH = 33;
  localparam int SCRATCHPAD_NUM_FILTER_BLOCKS_PER_MEGABLOCK = 1;
  localparam int SCRATCHPAD_NUM_BIAS_SCALE_BLOCKS_PER_MEGABLOCK = 1;
  localparam int MAX_XBAR_INPUT_INTERFACES = 5;
  localparam int MAX_XBAR_OUTPUT_INTERFACES = 5;
  localparam int AUX_XBAR_INPUT_COUNTER_WIDTH = 24;
  localparam int AUX_XBAR_OUTPUT_COUNTER_WIDTH = 24;
  localparam bit ENABLE_ACTIVATION = 1;
  localparam bit ENABLE_DEPTHWISE = 0;
  localparam int XBAR_ID_DEPTHWISE = -1;
  localparam int CONFIG_ID_DEPTHWISE = -1;
  localparam bit ENABLE_DEPTHWISE_FILTER_BIAS = 0;
  localparam int XBAR_ID_DEPTHWISE_FILTER_BIAS = -1;
  localparam int CONFIG_ID_DEPTHWISE_FILTER_BIAS = -1;
  localparam bit ENABLE_POOL = 1;
  localparam bit ENABLE_SOFTMAX = 1;
  localparam int XBAR_ID_SOFTMAX = 3;
  localparam int XBAR_ID_POOL = 2;
  localparam int XBAR_ID_ACTIVATION = 1;
  localparam int XBAR_ID_XBAR_OUT_PORT = 0;
  localparam int XBAR_ID_PE_ARRAY = 0;
  localparam int NUMBER_OF_KERNELS = 3;
  localparam int AUX_MODULE_SELECT_ID_WIDTH = 4;
  localparam bit XBAR_KERNEL_BYPASS_FEATURE_ENABLE = 0;
  localparam bit AUX_KERNEL_BYPASSABLE [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0};
  localparam int AUX_XBAR_MUX_OUTPUT_PIPELINE_STAGES [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0};
  localparam int AUX_XBAR_NONSTALLABLE_OUTPUT_PIPELINE_STAGES [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0};
  localparam int AUX_XBAR_OUTPUT_BP_FIFO_ENABLE [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0};
  localparam int AUX_XBAR_OUTPUT_BP_FIFO_DEPTH [16:0] = '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0,default : 0};
  localparam int AUX_XBAR_OUTPUT_WIDTH = 64;
  localparam int AUX_OUTPUT_DATA_WIDTHS [16:0] = '{0:64,1:64,2:64,3:64,4:64,5:64,6:64,7:64,8:64,9:64,10:64,11:64,12:64,13:64,14:64,15:64,16:64,default : 0};
  localparam int AUX_INPUT_DATA_WIDTHS [16:0] = '{0:64,1:64,2:64,3:64,4:64,5:64,6:64,7:64,8:64,9:64,10:64,11:64,12:64,13:64,14:64,15:64,16:64,default : 0};
  localparam int AUX_MAX_DATABUS_WIDTH = 64;
  localparam int XBAR_KERNEL_CV_FEATURE_ENABLE = 1;
  localparam int AUX_KERNEL_CONNECTIVITY_VECTOR [16:0] [16:0] = '{0: '{0:1,1:1,2:1,3:1,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},1: '{0:1,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},2: '{0:1,1:1,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},3: '{0:1,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},4: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},5: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},6: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},7: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},8: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},9: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},10: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},11: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},12: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},13: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},14: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},15: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0},16: '{0:0,1:0,2:0,3:0,4:0,5:0,6:0,7:0,8:0,9:0,10:0,11:0,12:0,13:0,14:0,15:0,16:0}};
  localparam int ACTIVATION_K_VECTOR = 4;
  localparam bit ACTIVATION_ENABLE_DSP_MULT = 0;
  localparam bit ACTIVATION_ENABLE_DSP_CONV = 0;
  localparam int ACTIVATION_GROUP_DELAY = 1;
  localparam int ACTIVATION_TYPE = 1;
  localparam int ACTIVATION_PARAM_CACHE_DEPTH = 2048;
  localparam int POOL_K_VECTOR = 4;
  localparam int POOL_GROUP_DELAY = 1;
  localparam int POOL_TYPE = 0;
  localparam int POOL_CONFIG_ID_WIDTH = 1;
  localparam int POOL_MAX_WINDOW_HEIGHT = 3;
  localparam int POOL_MAX_WINDOW_WIDTH = 3;
  localparam int POOL_MAX_STRIDE_VERTICAL = 4;
  localparam int POOL_MAX_STRIDE_HORIZONTAL = 4;
  localparam int POOL_PIPELINE_REG_NUM = 1;
  localparam int DEPTHWISE_K_VECTOR = 0;
  localparam int DEPTHWISE_GROUP_DELAY = 1;
  localparam int DEPTHWISE_TYPE = 0;
  localparam int DEPTHWISE_CONFIG_ID_WIDTH = 1;
  localparam int DEPTHWISE_MAX_WINDOW_HEIGHT = 3;
  localparam int DEPTHWISE_MAX_WINDOW_WIDTH = 3;
  localparam int DEPTHWISE_MAX_STRIDE_VERTICAL = 4;
  localparam int DEPTHWISE_MAX_STRIDE_HORIZONTAL = 4;
  localparam int DEPTHWISE_PIPELINE_REG_NUM = 1;
  localparam int DEPTHWISE_MAX_DILATION_VERTICAL = 1;
  localparam int DEPTHWISE_MAX_DILATION_HORIZONTAL = 1;
  localparam int DEPTHWISE_VECTOR_FEATURE_WIDTH = 16;
  localparam int DEPTHWISE_VECTOR_FILTER_WIDTH = 16;
  localparam int DEPTHWISE_VECTOR_BIAS_WIDTH = 32;
  localparam int DEPTHWISE_VECTOR_DOT_SIZE = 10;
  localparam int SOFTMAX_K_VECTOR = 1;
  localparam int SOFTMAX_GROUP_DELAY = 1;
  localparam int SOFTMAX_CONFIG_ID_WIDTH = 8;
  localparam int SOFTMAX_MAX_NUM_CHANNELS = 16;
  localparam int AUX_MAX_TILE_HEIGHT = 128;
  localparam int AUX_MAX_TILE_WIDTH = 128;
  localparam int AUX_MAX_TILE_CHANNELS = 8192;
  localparam bit LAYOUT_TRANSFORM_ENABLE_IN_BIAS_SCALE = 0;
  localparam int LAYOUT_TRANSFORM_ENABLE = 0;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_ENABLE = 1;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_CHANNELS = 1;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_BUS_WIDTH = 128;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_ELEMENT_WIDTH = 16;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_PIXEL_FIFO_DEPTH = 16;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_CONV_MODE = 0;
  localparam int LIGHTWEIGHT_LAYOUT_TRANSFORM_BIAS_SCALE_ENABLE = 0;
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_CHANNELS = 3;
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_HEIGHT = 28;
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_WIDTH = 28;
  localparam int LAYOUT_TRANSFORM_MAX_FEATURE_DEPTH = 1;
  localparam int LAYOUT_TRANSFORM_MAX_STRIDE_WIDTH = 2;
  localparam int LAYOUT_TRANSFORM_MAX_STRIDE_HEIGHT = 2;
  localparam int LAYOUT_TRANSFORM_MAX_STRIDE_DEPTH = 1;
  localparam int LAYOUT_TRANSFORM_MAX_PAD_FRONT = 1;
  localparam int LAYOUT_TRANSFORM_MAX_PAD_LEFT = 2;
  localparam int LAYOUT_TRANSFORM_MAX_PAD_TOP = 2;
  localparam int LAYOUT_TRANSFORM_MAX_FILTER_HEIGHT = 2;
  localparam int LAYOUT_TRANSFORM_MAX_FILTER_WIDTH = 2;
  localparam int LAYOUT_TRANSFORM_MAX_FILTER_DEPTH = 1;
  localparam int LAYOUT_TRANSFORM_MAX_DILATION_WIDTH = 2;
  localparam int LAYOUT_TRANSFORM_MAX_DILATION_HEIGHT = 2;
  localparam int LAYOUT_TRANSFORM_MAX_DILATION_DEPTH = 1;
  localparam int LAYOUT_TRANSFORM_READER_BYTES = 16;
  localparam int LAYOUT_TRANSFORM_CONV_MODE = 0;
  localparam int ENABLE_OUTPUT_STREAMER = 1;
  localparam int AXI_OSTREAM_DATA_WIDTH = 128;
  localparam int AXI_OSTREAM_ID_WIDTH = 8;
  localparam int AXI_OSTREAM_DEST_WIDTH = 8;
  localparam int AXI_OSTREAM_FIFO_DEPTH = 128;
  localparam int DISABLE_DDR = 1;
`endif // DLA_DMA_PARAM_SVH
