// Copyright 2015-2020 Altera Corporation.
//
// This software and the related documents are Altera copyrighted materials,
// and your use of them is governed by the express license under which they
// were provided to you ("License"). Unless the License provides otherwise,
// you may not use, modify, copy, publish, distribute, disclose or transmit
// this software or the related documents without Altera's prior written
// permission.
//
// This software and the related documents are provided as is, with no express
// or implied warranties, other than those that are expressly stated in the
// License.

// --- dla_top_derived_params.sv -----------------------------------------------
// This file contains derived parameters that are calculated based on the
// top-level parameters to dla_top.
// -----------------------------------------------------------------------------

localparam int BYTE_WIDTH = 8;
localparam int FP16_WIDTH = 16;

localparam int FILTER_READER_WIDTH = FILTER_READER_DATA_BYTES*BYTE_WIDTH;
localparam int FEATURE_READER_WIDTH = FEATURE_READER_DATA_BYTES*BYTE_WIDTH;
localparam int FEATURE_WRITER_WIDTH = FEATURE_WRITER_DATA_BYTES*BYTE_WIDTH;
localparam int CONFIG_READER_WIDTH = CONFIG_READER_DATA_BYTES*BYTE_WIDTH;
localparam int CONFIG_WIDTH = CONFIG_DATA_BYTES*BYTE_WIDTH;


localparam dla_pe_array_pkg::pe_array_arch_t PE_ARRAY_ARCH = dla_pe_array_pkg::pe_array_arch_t'(PE_ARRAY_PARAM_BITS);

localparam int PE_ARRAY_LANE_DATA_WIDTH = PE_ARRAY_ARCH.NUM_RESULTS_PER_CYCLE * FP16_WIDTH;

// The input_feeder accepts input data that is sized to be stored in the stream
// buffer and then sent to the PE array without having to be resized further.
// Therefore, the input width of the input_feeder depends on the PE array block
// size (C_VECTOR).
localparam int INPUT_FEEDER_LANE_DATA_WIDTH = PE_ARRAY_ARCH.DOT_SIZE * FP16_WIDTH;

`include "dla_pe_array_constants.svh"

localparam int SCRATCHPAD_NUM_PE_PORTS = PE_ARRAY_ARCH.NUM_PES * PE_ARRAY_ARCH.NUM_FILTERS;
localparam int SCRATCHPAD_NUM_READ_BRANCH_PIPELINE = 1;
localparam int SCRATCHPAD_NUM_READ_PIPELINE_CYCLE = 1;

localparam int PE_ARRAY_EXIT_FIFO_ALMOST_FULL_CUTOFF = get_total_pe_array_latency(PE_ARRAY_ARCH) + SCRATCHPAD_ARCH_INFO.READ_TO_OUTPUT_DELAY;

localparam int SCRATCHPAD_MEM_ID_WIDTH =
  dla_filter_bias_scale_scratchpad_pkg::calc_mem_id_width(
    .NUM_PE_PORTS(SCRATCHPAD_NUM_PE_PORTS),
    .NUM_FILTER_PORTS(SCRATCHPAD_NUM_FILTER_PORTS),
    .NUM_BIAS_SCALE_PORTS(SCRATCHPAD_NUM_BIAS_SCALE_PORTS));
localparam int SCRATCHPAD_MEM_ADDR_WIDTH =
  dla_filter_bias_scale_scratchpad_pkg::calc_mem_addr_width(
    .FILTER_DEPTH(SCRATCHPAD_FILTER_DEPTH),
    .BIAS_SCALE_DEPTH(SCRATCHPAD_BIAS_SCALE_DEPTH));
localparam int SCRATCHPAD_FILTER_BASE_ADDR_WIDTH =
  dla_filter_bias_scale_scratchpad_pkg::calc_filter_base_addr_width(
    .FILTER_DEPTH(SCRATCHPAD_FILTER_DEPTH));
localparam int SCRATCHPAD_BIAS_SCALE_BASE_ADDR_WIDTH =
  dla_filter_bias_scale_scratchpad_pkg::calc_bias_scale_base_addr_width(
    .BIAS_SCALE_DEPTH(SCRATCHPAD_BIAS_SCALE_DEPTH));

localparam device_family_t DEVICE_ENUM = PE_ARRAY_ARCH.DEVICE;

// Parameter checking.
initial begin
  if (DEVICE_ENUM == -1) begin
    $fatal(1, "DEVICE was not set to a valid value");
  end

  if (PE_ARRAY_ARCH.DOT_MODE == -1) begin
    $fatal(1, "PE_ARRAY_DOT_MODE was not set to a valid value");
  end

  if (PE_ARRAY_ARCH.CONVERT_MODE == -1) begin
    $fatal(1, "PE_ARRAY_CONVERT_MODE was not set to a valid value");
  end

  if (PE_ARRAY_ARCH.ACCUM_MODE == -1) begin
    $fatal(1, "PE_ARRAY_ACCUM_MODE was not set to a valid value");
  end
end

localparam dla_aux_depthwise_pkg::vector_dot_arch_t AUX_DEPTHWISE_VECTOR_ARCH = '{
  FEATURE_WIDTH :  DEPTHWISE_VECTOR_FEATURE_WIDTH,
  FILTER_WIDTH  :  DEPTHWISE_VECTOR_FILTER_WIDTH,
  BIAS_WIDTH    :  DEPTHWISE_VECTOR_BIAS_WIDTH,
  DOT_SIZE      :  DEPTHWISE_VECTOR_DOT_SIZE,
  DEVICE        :  DEVICE_ENUM
};

localparam dla_aux_depthwise_pkg::vector_dot_arch_info_t DEPTHWISE_VECTOR_ARCH_INFO = dla_aux_depthwise_pkg::get_arch_info(AUX_DEPTHWISE_VECTOR_ARCH);

localparam dla_filter_bias_scale_scratchpad_pkg::filter_bias_scale_scratchpad_arch_t SCRATCHPAD_ARCH = '{
  DEVICE: DEVICE_ENUM,
  NUM_PE_PORTS: SCRATCHPAD_NUM_PE_PORTS,
  FILTER_DEPTH: SCRATCHPAD_FILTER_DEPTH,
  BIAS_SCALE_DEPTH: SCRATCHPAD_BIAS_SCALE_DEPTH,
  NUM_FILTER_PORTS: SCRATCHPAD_NUM_FILTER_PORTS,
  NUM_BIAS_SCALE_PORTS: SCRATCHPAD_NUM_BIAS_SCALE_PORTS,
  NUM_READ_PIPELINE_MEM: PE_ARRAY_ARCH.NUM_FILTERS,
  NUM_WRITE_PIPELINE_MEM: PE_ARRAY_ARCH.NUM_FILTERS,
  NUM_READ_BRANCH_PIPELINE: SCRATCHPAD_NUM_READ_BRANCH_PIPELINE,
  NUM_READ_PIPELINE_CYCLE: SCRATCHPAD_NUM_READ_PIPELINE_CYCLE,
  ENABLE_SCALE: PE_ARRAY_ARCH.ENABLE_SCALE,
  ENABLE_DDRFREE_FBS: PE_ARRAY_ARCH.ENABLE_DDRFREE_FBS,
  BLOCK_SIZE: PE_ARRAY_ARCH.DOT_SIZE,
  FILTER_WIDTH: PE_ARRAY_ARCH.FILTER_WIDTH,
  FILTER_EXPONENT_WIDTH: PE_ARRAY_ARCH.FILTER_EXPONENT_WIDTH,
  BIAS_WIDTH: BIAS_WIDTH,
  SCALE_WIDTH: SCALE_WIDTH,

  MEGABLOCK_WIDTH: SCRATCHPAD_MEGABLOCK_WIDTH,
  NUM_FILTER_BLOCKS_PER_MEGABLOCK: SCRATCHPAD_NUM_FILTER_BLOCKS_PER_MEGABLOCK,
  NUM_BIAS_SCALE_BLOCKS_PER_MEGABLOCK: SCRATCHPAD_NUM_BIAS_SCALE_BLOCKS_PER_MEGABLOCK
};

localparam dla_filter_bias_scale_scratchpad_pkg::filter_bias_scale_scratchpad_arch_info_t SCRATCHPAD_ARCH_INFO =
  dla_filter_bias_scale_scratchpad_pkg::get_arch_info(SCRATCHPAD_ARCH);


localparam int SCRATCHPAD_LATENCY = SCRATCHPAD_ARCH_INFO.READ_TO_OUTPUT_DELAY;

localparam int PE_ARRAY_VALID_LATENCY = SCRATCHPAD_LATENCY;

localparam int PE_ARRAY_FLUSH_LATENCY = 0; // Deprecated

localparam int PE_ARRAY_RESULT_ID_LATENCY = 0; // Deprecated

localparam dla_sequencer_pkg::sequencer_arch_t SEQUENCER_ARCH = '{
  ELTWISE_MULT_CMD_WIDTH: PE_ARRAY_ARCH.ELTWISE_MULT_CMD_WIDTH,
  RESULT_ID_WIDTH: PE_ARRAY_ARCH.RESULT_ID_WIDTH,

  SCRATCHPAD_MEM_ID_WIDTH: SCRATCHPAD_MEM_ID_WIDTH,
  SCRATCHPAD_MEM_ADDR_WIDTH: SCRATCHPAD_MEM_ADDR_WIDTH,
  SCRATCHPAD_FILTER_BASE_ADDR_WIDTH: SCRATCHPAD_FILTER_BASE_ADDR_WIDTH,
  SCRATCHPAD_BIAS_SCALE_BASE_ADDR_WIDTH: SCRATCHPAD_BIAS_SCALE_BASE_ADDR_WIDTH,

  NUM_BIAS_ID: divceil(SCRATCHPAD_NUM_PE_PORTS, SCRATCHPAD_NUM_BIAS_SCALE_PORTS),
  NUM_FILTER_ID: divceil(SCRATCHPAD_NUM_PE_PORTS, SCRATCHPAD_NUM_FILTER_PORTS),
  FILTER_CACHE_DEPTH: SCRATCHPAD_FILTER_DEPTH,
  BIAS_CACHE_DEPTH: SCRATCHPAD_BIAS_SCALE_DEPTH,

  NUM_RESULT_ID: PE_ARRAY_ARCH.NUM_RESULT_ID,
  NUM_INTERLEAVED_FEATURES: PE_ARRAY_ARCH.NUM_INTERLEAVED_FEATURES,
  NUM_INTERLEAVED_FILTERS: PE_ARRAY_ARCH.NUM_INTERLEAVED_FILTERS,

  PE_ARRAY_VALID_LATENCY: PE_ARRAY_VALID_LATENCY,
  PE_ARRAY_FLUSH_LATENCY: PE_ARRAY_FLUSH_LATENCY,
  PE_ARRAY_RESULT_ID_LATENCY: PE_ARRAY_RESULT_ID_LATENCY,

  ENABLE_DDRFREE_FBS: PE_ARRAY_ARCH.ENABLE_DDRFREE_FBS,

  DEVICE: DEVICE_ENUM
};

localparam dla_input_feeder_pkg::input_feeder_arch_t INPUT_FEEDER_ARCH = '{
  STREAM_BUFFER_DEPTH: STREAM_BUFFER_DEPTH,
  CONFIG_WIDTH: CONFIG_WIDTH,

  C_VECTOR: PE_ARRAY_ARCH.DOT_SIZE,
  FEATURE_WIDTH: PE_ARRAY_ARCH.FEATURE_WIDTH,
  FEATURE_EXPONENT_WIDTH: PE_ARRAY_ARCH.FEATURE_EXPONENT_WIDTH,
  FEATURE_EXPONENT_BIAS: PE_ARRAY_ARCH.FEATURE_EXPONENT_BIAS,

  KVEC_OVER_CVEC: KVEC_OVER_CVEC,
  FILTER_ADDR_WIDTH: $clog2(SCRATCHPAD_FILTER_DEPTH),
  BIAS_ADDR_WIDTH: $clog2(SCRATCHPAD_BIAS_SCALE_DEPTH),

  NUM_INTERLEAVED_FEATURES: PE_ARRAY_ARCH.NUM_INTERLEAVED_FEATURES,
  NUM_INTERLEAVED_FILTERS: PE_ARRAY_ARCH.NUM_INTERLEAVED_FILTERS,

  NUM_LANES: PE_ARRAY_ARCH.NUM_LANES,
  NUM_FEATURES: PE_ARRAY_ARCH.NUM_FEATURES,
  FEATURE_READER_WIDTH: FEATURE_READER_WIDTH,
  GROUP_DELAY: PE_ARRAY_ARCH.GROUP_DELAY,

  ENABLE_DDRFREE_FBS: PE_ARRAY_ARCH.ENABLE_DDRFREE_FBS,
  ENABLE_MIXED_PRECISION: ENABLE_MIXED_PRECISION,
  DEVICE: DEVICE_ENUM
};

localparam dla_exit_fifo_pkg::exit_fifo_arch_t EXIT_FIFO_ARCH = '{
  NUM_LANES: PE_ARRAY_ARCH.NUM_LANES,
  NUM_RESULTS_PER_CYCLE: PE_ARRAY_ARCH.NUM_RESULTS_PER_CYCLE,
  NUM_FEATURES: PE_ARRAY_ARCH.NUM_FEATURES,

  FIFO_DEPTH: PE_ARRAY_EXIT_FIFO_DEPTH,
  FIFO_ALMOST_FULL_CUTOFF: PE_ARRAY_EXIT_FIFO_ALMOST_FULL_CUTOFF,
  GROUP_DELAY: PE_ARRAY_ARCH.GROUP_DELAY
};

localparam int LT_ELEMENT_WIDTH = LAYOUT_TRANSFORM_CONV_MODE == U8_TO_F16 ? 8 : 16;
localparam dla_lt_pkg::lt_arch_t LT_ARCH = '{
  ENABLE_LT: LAYOUT_TRANSFORM_ENABLE,
  ENABLE_IN_BIAS_SCALE: LAYOUT_TRANSFORM_ENABLE_IN_BIAS_SCALE,
  KEEP_SINGLE_CONFIG: ENABLE_ON_CHIP_PARAMETERS,
  DATA_ELEMENT_WIDTH: LT_ELEMENT_WIDTH,
  CNT_BITS: 20,
  CONV_MODE: dla_lt_pkg::convert_mode_t'(LAYOUT_TRANSFORM_CONV_MODE),
  DDR_BYTES: LAYOUT_TRANSFORM_READER_BYTES,
  CONFIG_BYTES: CONFIG_DATA_BYTES,
  MAX_CHANNELS: LAYOUT_TRANSFORM_MAX_FEATURE_CHANNELS,
  MAX_FEATURE_HEIGHT: LAYOUT_TRANSFORM_MAX_FEATURE_HEIGHT,
  MAX_FEATURE_WIDTH: LAYOUT_TRANSFORM_MAX_FEATURE_WIDTH,
  MAX_FEATURE_DEPTH: LAYOUT_TRANSFORM_MAX_FEATURE_DEPTH,
  MAX_STRIDE_HEIGHT: LAYOUT_TRANSFORM_MAX_STRIDE_HEIGHT,
  MAX_STRIDE_WIDTH: LAYOUT_TRANSFORM_MAX_STRIDE_WIDTH,
  MAX_STRIDE_DEPTH: LAYOUT_TRANSFORM_MAX_STRIDE_DEPTH,
  CVEC: PE_ARRAY_ARCH.DOT_SIZE,
  MAX_PAD_FRONT: LAYOUT_TRANSFORM_MAX_PAD_FRONT,
  MAX_PAD_LEFT: LAYOUT_TRANSFORM_MAX_PAD_LEFT,
  MAX_PAD_TOP: LAYOUT_TRANSFORM_MAX_PAD_TOP,
  MAX_FILTER_HEIGHT: LAYOUT_TRANSFORM_MAX_FILTER_HEIGHT,
  MAX_FILTER_WIDTH: LAYOUT_TRANSFORM_MAX_FILTER_WIDTH,
  MAX_FILTER_DEPTH: LAYOUT_TRANSFORM_MAX_FILTER_DEPTH,
  MAX_DILATION_HEIGHT: LAYOUT_TRANSFORM_MAX_DILATION_HEIGHT,
  MAX_DILATION_WIDTH: LAYOUT_TRANSFORM_MAX_DILATION_WIDTH,
  MAX_DILATION_DEPTH: LAYOUT_TRANSFORM_MAX_DILATION_DEPTH,
  DEVICE: DEVICE_ENUM
};

localparam dla_lw_lt_pkg::lw_lt_arch_t LW_LT_ARCH = '{
  LW_LT_ENABLED: LIGHTWEIGHT_LAYOUT_TRANSFORM_ENABLE,
  CONFIG_BYTES: CONFIG_DATA_BYTES,
  CVEC: PE_ARRAY_ARCH.DOT_SIZE,
  AXI_WIDTH: LIGHTWEIGHT_LAYOUT_TRANSFORM_BUS_WIDTH,
  CHANNELS: LIGHTWEIGHT_LAYOUT_TRANSFORM_CHANNELS,
  CONV_MODE: dla_lt_pkg::convert_mode_t'(LIGHTWEIGHT_LAYOUT_TRANSFORM_CONV_MODE),
  DEVICE: DEVICE_ENUM,
  ENABLE_IN_BIAS_SCALE: LIGHTWEIGHT_LAYOUT_TRANSFORM_BIAS_SCALE_ENABLE,
  PIXEL_EXIT_FIFO_DEPTH: LIGHTWEIGHT_LAYOUT_TRANSFORM_PIXEL_FIFO_DEPTH
};
